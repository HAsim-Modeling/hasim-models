`include "hasim_common.bsh"
`include "hasim_core.bsh"

module [HASIM_MODULE] mkChip();
    let core <- mkCore;
endmodule
