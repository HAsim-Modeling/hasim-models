`include "hasim_common.bsh"

module [HASIM_MODULE] mkMemory();
    return ?;
endmodule
