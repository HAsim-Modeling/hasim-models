`include "hasim_common.bsh"
`include "hasim_pipeline.bsh"

module [HASIM_MODULE] mkCore();
    let pipeline <- mkPipeline;
endmodule
