`include "asim/provides/hasim_common.bsh"
`include "asim/provides/hasim_pipeline.bsh"

module [HASIM_MODULE] mkCore();
    let pipeline <- mkPipeline;
endmodule
