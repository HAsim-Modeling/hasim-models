//
// Copyright (c) 2014, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//
// ******* Library Imports *******

import Vector::*;
import FIFO::*;

// ******* Application Imports *******

`include "awb/provides/soft_connections.bsh"
`include "awb/provides/common_services.bsh"
`include "awb/provides/fpga_components.bsh"


// ******* HAsim Imports *******

`include "awb/provides/hasim_common.bsh"
`include "awb/provides/hasim_model_services.bsh"
`include "awb/provides/hasim_modellib.bsh"

`include "awb/provides/funcp_base_types.bsh"
`include "awb/provides/funcp_memstate_base_types.bsh"
`include "awb/provides/funcp_interface.bsh"


// ******* Timing Model Imports *******

`include "awb/provides/memory_base_types.bsh"
`include "awb/provides/chip_base_types.bsh"
`include "awb/provides/hasim_cache_protocol.bsh"
`include "awb/provides/hasim_cache_algorithms.bsh"
`include "awb/provides/hasim_l2_cache_alg.bsh"
`include "awb/provides/hasim_miss_tracker.bsh"

// ******* Generated File Imports *******

`include "awb/dict/EVENTS_L2.bsh"


// ****** Local Definitions *******


typedef `L2_MISS_ID_SIZE L2_MISS_ID_SIZE;
typedef CACHE_MISS_INDEX#(L2_MISS_ID_SIZE) L2_MISS_ID;
typedef CACHE_MISS_TOKEN#(L2_MISS_ID_SIZE) L2_MISS_TOKEN;
typedef TExp#(L2_MISS_ID_SIZE) NUM_L2_MISS_IDS;

typedef enum
{
    L2_CC_REQ_WB,
    L2_CC_REQ_INVALIDATE
}
L2_CC_REQ deriving (Eq, Bits);


//
// L2_LOCAL_STATE --
//   L2 State to pass between pipeline stages.
//
typedef struct
{
    L2_MISS_TOKEN missTokToFree;

    Bool memQNotFull;
    Bool memQUsed;
    CACHE_PROTOCOL_MSG memQData;
    
    Bool writePortUsed;
    L2_CACHE_IDX writePortIdx;
    CACHE_ENTRY_STATE#(void) writePortData;
    
    Bool coreQNotFull;
    Bool coreQUsed;
    CACHE_PROTOCOL_MSG coreQData;

    Maybe#(CACHE_PROTOCOL_MSG) req;
}
L2_LOCAL_STATE deriving (Eq, Bits);

// initLocalState
//
// A fresh local state for the first stage.

function L2_LOCAL_STATE initLocalState();
    return 
        L2_LOCAL_STATE 
        { 
            missTokToFree: ?,
            memQNotFull: True,
            memQUsed: False,
            memQData: ?,
            coreQNotFull: True,
            coreQUsed: False,
            coreQData: ?,
            writePortUsed: False,
            writePortIdx: ?,
            writePortData: ?,
            req: tagged Invalid
        };
endfunction

//
// memQAvailable --
//   The memQ is available if it is notFull AND someone has
//   not already used it.
//
function Bool memQAvailable(L2_LOCAL_STATE local_state);
    return local_state.memQNotFull && !local_state.memQUsed;
endfunction


// mkL2Cache

// A model of an L2 Cache that is unpipelined.
// That is, writes to the cache occur in the same model cycle as hit checks.
// In a more realistic model a writeQ would track pending updates.
// Also there is no victim buffer.
//
// Note that the module itself is implemented as a pipeline, though the target
// model carries out all actions in one model cycle.

module [HASIM_MODULE] mkL2Cache#(String reqFromL1Name,
                                 String rspToL1Name,
                                 String reqToMemoryName,
                                 String rspFromMemoryName)
    // Interface:
    ();

    TIMEP_DEBUG_FILE_MULTIPLEXED#(MAX_NUM_CPUS) debugLog <- mkTIMEPDebugFile_Multiplexed("cache_l2_data.out");

    // ****** Submodels ******

    // The cache algorithm which determines hits, misses, and evictions.
    function Bool alwaysTrue(t_DUMMY d) = True;
    L2_CACHE_ALG#(MAX_NUM_CPUS, void) l2Alg <- mkL2CacheAlg(alwaysTrue);

    // Track the next Miss ID to give out.
    CACHE_MISS_TRACKER#(MAX_NUM_CPUS, L2_MISS_ID_SIZE) outstandingMisses <- mkCacheMissTracker();

    // A RAM To map our miss IDs into the original opaques, that we return to higher levels.
    MEMORY_IFC_MULTIPLEXED#(MAX_NUM_CPUS, L2_MISS_ID,
                            Tuple2#(L2_MISS_TOKEN, L2_CACHE_IDX)) opaquesPool <-
        mkMemory_Multiplexed(mkBRAM);

    // ****** Ports ******

    // Queues to/from core hierarchy.
    PORT_STALL_RECV_MULTIPLEXED#(MAX_NUM_CPUS, CACHE_PROTOCOL_MSG) reqFromCore <-
        mkPortStallRecv_Multiplexed(reqFromL1Name);
    PORT_STALL_SEND_MULTIPLEXED#(MAX_NUM_CPUS, CACHE_PROTOCOL_MSG) rspToCore <-
        mkPortStallSend_Multiplexed(rspToL1Name);
    
    // Queues to/from coherence engine.
    PORT_STALL_SEND_MULTIPLEXED#(MAX_NUM_CPUS, MEMORY_REQ) reqToUncore <-
        mkPortStallSend_Multiplexed(reqToMemoryName);
    
    PORT_STALL_RECV_MULTIPLEXED#(MAX_NUM_CPUS, MEMORY_RSP) rspFromUncore <-
        mkPortStallRecv_Multiplexed(rspFromMemoryName);
    
    Vector#(4, INSTANCE_CONTROL_IN#(MAX_NUM_CPUS))  inctrls = newVector();
    Vector#(4, INSTANCE_CONTROL_OUT#(MAX_NUM_CPUS)) outctrls = newVector();
    
    inctrls[0]  = reqFromCore.ctrl.in;
    inctrls[1]  = rspToCore.ctrl.in;
    inctrls[2]  = reqToUncore.ctrl.in;
    inctrls[3]  = rspFromUncore.ctrl.in;

    outctrls[0] = reqFromCore.ctrl.out;
    outctrls[1] = rspToCore.ctrl.out;
    outctrls[2] = reqToUncore.ctrl.out;
    outctrls[3] = rspFromUncore.ctrl.out;

    LOCAL_CONTROLLER#(MAX_NUM_CPUS) localCtrl <- mkNamedLocalController("L2 Cache", inctrls, outctrls);

    STAGE_CONTROLLER#(MAX_NUM_CPUS, L2_LOCAL_STATE) stage2Ctrl <- mkBufferedStageController();
    STAGE_CONTROLLER#(MAX_NUM_CPUS, L2_LOCAL_STATE) stage3Ctrl <- mkBufferedStageController();
    STAGE_CONTROLLER#(MAX_NUM_CPUS, L2_LOCAL_STATE) stage4Ctrl <- mkBufferedStageController();
    STAGE_CONTROLLER#(MAX_NUM_CPUS, Tuple3#(L2_LOCAL_STATE,
                                            Maybe#(CACHE_PROTOCOL_MSG),
                                            L2_CACHE_IDX)) stage5Ctrl <-
        mkStageController();

    Reg#(Maybe#(Tuple4#(CPU_INSTANCE_ID,
                        CACHE_PROTOCOL_MSG,
                        L2_CACHE_LOOKUP_RSP#(void),
                        L2_LOCAL_STATE))) stage4Stall <- mkReg(tagged Invalid);


    // ****** Stats ******

    STAT_VECTOR#(MAX_NUM_CPUS) statReadHit <-
        mkStatCounter_Multiplexed(statName("MODEL_L2_READ_HIT",
                                           "L2 Read Hits"));
    STAT_VECTOR#(MAX_NUM_CPUS) statReadMiss <-
        mkStatCounter_Multiplexed(statName("MODEL_L2_READ_MISS",
                                           "L2 Read Misses"));
    STAT_VECTOR#(MAX_NUM_CPUS) statReadRetry <-
        mkStatCounter_Multiplexed(statName("MODEL_L2_READ_RETRY",
                                           "L2 Read Retries"));
    STAT_VECTOR#(MAX_NUM_CPUS) statWriteHit <-
        mkStatCounter_Multiplexed(statName("MODEL_L2_WRITE_HIT",
                                           "L2 Write Hits"));
    STAT_VECTOR#(MAX_NUM_CPUS) statWriteRetry <-
        mkStatCounter_Multiplexed(statName("MODEL_L2_WRITE_RETRY",
                                           "L2 Write Retries"));
    STAT_VECTOR#(MAX_NUM_CPUS) statFillRetry <-
        mkStatCounter_Multiplexed(statName("MODEL_L2_FILL_RETRY",
                                           "L2 Fill Retries"));

    EVENT_RECORDER_MULTIPLEXED#(MAX_NUM_CPUS) eventHit  <- mkEventRecorder_Multiplexed(`EVENTS_L2_HIT);
    EVENT_RECORDER_MULTIPLEXED#(MAX_NUM_CPUS) eventMiss <- mkEventRecorder_Multiplexed(`EVENTS_L2_MISS);
    EVENT_RECORDER_MULTIPLEXED#(MAX_NUM_CPUS) eventFill <- mkEventRecorder_Multiplexed(`EVENTS_L2_FILL);

    // ****** Assertions ******

    let assertReqOk <- mkAssertionSimOnly("l2-cache-controller-unpipelined.bsv: Unexpected request kind",
                                          ASSERT_ERROR);
    let assertRspOk <- mkAssertionSimOnly("l2-cache-controller-unpipelined.bsv: Unexpected response kind",
                                          ASSERT_ERROR);


    //
    // Stage 1 --
    //   Consume responses from memory.
    //
    (* conservative_implicit_conditions *)
    rule stage1_fill (True);
        // Start a new model cycle
        let cpu_iid <- localCtrl.startModelCycle();
        debugLog.nextModelCycle(cpu_iid);

        // Make a conglomeration of local information to pass from stage to stage.
        let local_state = initLocalState();

        // Check if the CC engine has room for any new requests.
        let can_enq_uncore_req <- reqToUncore.canEnq(cpu_iid);
        let can_enq_core_rsp <- rspToCore.canEnq(cpu_iid);
        local_state.memQNotFull = can_enq_uncore_req;
        local_state.coreQNotFull = can_enq_core_rsp;
        
        // Now check for responses from the cache coherence engine.
        let m_uncore_rsp <- rspFromUncore.receive(cpu_iid);

        Bool read_opaques = False;

        //
        // Have a response from memory?
        //
        if (m_uncore_rsp matches tagged Valid .mem_rsp)
        begin
            let rsp = cacheMsgFromMemRsp(mem_rsp);

            assertRspOk(cacheMsg_IsRspLoad(rsp));

            // Yes.  Can it be sent up toward the core?
            if (local_state.coreQNotFull)
            begin
                // Yes.  Consume the response.
                let fill = rsp;

                // We want to use the cache write port.
                // Since we're the highest priority we don't have to check if
                // someone else has it. Just record that we're using it so
                // no one else will.
                local_state.writePortUsed = True;
                local_state.writePortData = initCacheEntryState(fill.linePAddr,
                                                                False,
                                                                ?);

                // Get the Miss ID.
                L2_MISS_TOKEN miss_tok = fromMemOpaque(fill.opaque);

                // Free the token in the next stage, in case we had to retry.
                local_state.missTokToFree = miss_tok;

                // Return the fill to higher levels.
                debugLog.record_next_cycle(cpu_iid, $format("1: MEM RSP: %0d, LINE: 0x%h", miss_tok.index, fill.linePAddr));

                // Read the meta-data from the fill request
                opaquesPool.readReq(cpu_iid, missTokIndex(miss_tok));

                // Only respond to loads.
                if (missTokIsLoad(miss_tok))
                begin
                    local_state.coreQUsed = True;
                    local_state.coreQData = fill;
                end
            end
            else
            begin
                // Can't consume the response because there is no space to
                // forward it. 
                L2_MISS_TOKEN miss_tok = fromMemOpaque(rsp.opaque);
                debugLog.record_next_cycle(cpu_iid, $format("1: MEM RSP RETRY: %0d, LINE: 0x%h", miss_tok.index, rsp.linePAddr));
            end
        end
        else
        begin
            // There's no response from the below.
            debugLog.record_next_cycle(cpu_iid, $format("1: NO MEM RSP"));
        end

        stage2Ctrl.ready(cpu_iid, local_state);
    endrule


    //
    // stage2_victimIdx --
    //   Learn the index of the victim and check the victim line's current state.
    //
    rule stage2_victimIdx (True);
        match {.cpu_iid, .local_state} <- stage2Ctrl.nextReadyInstance();

        if (local_state.writePortUsed)
        begin
            match {.prev_opaque, .fill_idx} <- opaquesPool.readRsp(cpu_iid);

            // Record the cache fill index
            local_state.writePortIdx = fill_idx;

            //
            // Restore the opaque to the context that sent the request to this
            // cache.  This cache modified only the bits required for a local
            // miss token.  Merge the unmodified bits (still in the opaque)
            // and the preserved, overwritten bits (stored in opaquesPool).
            //
            if (local_state.coreQUsed)
            begin
                local_state.coreQData.opaque = updateMemOpaque(local_state.coreQData.opaque,
                                                               prev_opaque);
            end

            // Does the current entry that will be evicted need writeback?
            l2Alg.lookupByIndexReq(cpu_iid, fill_idx);
        end

        stage3Ctrl.ready(cpu_iid, local_state);
    endrule


    //
    // stage3_evictAndCPUReq --
    //   Finish fill evictions and request lookups for any load/stores.
    //
    rule stage3_evictAndCPUReq (True);
        match {.cpu_iid, .local_state} <- stage3Ctrl.nextReadyInstance();

        // See if we started an eviction in the previous stage.
        if (local_state.writePortUsed)
        begin
            let m_evict <- l2Alg.lookupByIndexRsp(cpu_iid);

            // If our fill evicted a dirty line we must write it back.
            if (m_evict matches tagged Valid .state &&&
                state.dirty)
            begin
                // Is there any room in the memQ?
                if (memQAvailable(local_state))
                begin
                    debugLog.record(cpu_iid, $format("2: DIRTY EVICTION: 0x%h", state.linePAddr));

                    // Record that we're using the memQ.
                    local_state.memQUsed = True;
                    local_state.memQData = cacheMsg_ReqStore(state.linePAddr, ?);
                    outstandingMisses.free(cpu_iid, local_state.missTokToFree);
                
                    // Acknowledge the fill.
                    rspFromUncore.doDeq(cpu_iid);
                end
                else
                begin
                    // The queue is full, so retry the fill next cycle. No dequeue.
                    rspFromUncore.noDeq(cpu_iid);
                    
                    debugLog.record(cpu_iid, $format("2: DIRTY EVICTION RETRY: 0x%h", state.linePAddr));

                    // Yield the writePort and rspPort to lower-priority users.
                    // The fill update will not happen this model cycle.
                    // Don't free the token.
                    local_state.writePortUsed = False;
                    local_state.coreQUsed = False;
                end
            end
            else
            begin
                // We finished the fill succesfully and no writeback is needed.
                // Dequeue the fill and free the miss.
                debugLog.record(cpu_iid, $format("2: CLEAN EVICTION"));
                outstandingMisses.free(cpu_iid, local_state.missTokToFree);
                rspFromUncore.doDeq(cpu_iid);
            end

            // Note that the actual cache update will be done later, so that
            // any lookups this model cycle don't see it accidentally.
        end
        else
        begin
            // No fill received
            rspFromUncore.noDeq(cpu_iid);
        end

        if (local_state.writePortUsed)
        begin
            eventFill.recordEvent(cpu_iid,
                                  tagged Valid resize({ local_state.writePortData.linePAddr, 1'b0 }));
        end
        else
        begin
            eventFill.recordEvent(cpu_iid, tagged Invalid);
        end


        // Now read the request port from the L1.
        let m_core_req <- reqFromCore.receive(cpu_iid);

        // Deal with any load/store requests.
        if (m_core_req matches tagged Valid .req)
        begin
            assertReqOk(cacheMsg_IsReqLoad(req) || cacheMsg_IsReqStore(req));

            // See if the cache algorithm hit or missed.
            l2Alg.lookupByAddrReq(cpu_iid,
                                  req.linePAddr,
                                  True,
                                  local_state.coreQUsed);
            debugLog.record(cpu_iid, $format("2: REQ: LINE: 0x%h", req.linePAddr));

            // Finish the request in the next stage.
            local_state.req = tagged Valid req;
        end
        else
        begin
            debugLog.record(cpu_iid, $format("2: NO REQ"));
        end
        
        // Pass our information to the next stage.
        stage4Ctrl.ready(cpu_iid, local_state);
    endrule
    
    
    //
    // stage4_cpuRspStoreReq --
    //   Finish up any load/stores to see if they hit or miss.
    //   Begin handling any store requests.
    //    
    rule stage4_cpuRspCCReq (!isValid(stage4Stall));
        // Get the local state from the previous stage.
        match {.cpu_iid, .local_state} <- stage4Ctrl.nextReadyInstance();

        // See if we need to finish any cpu responses.
        if (local_state.req matches tagged Valid .req)
        begin
            // Get the lookup response.
            let entry <- l2Alg.lookupByAddrRsp(cpu_iid);
            stage4Stall <= tagged Valid tuple4(cpu_iid, req, entry, local_state);
        end
        else
        begin
            // No request.  Propogate the bubble.
            reqFromCore.noDeq(cpu_iid);
            eventHit.recordEvent(cpu_iid, tagged Invalid);
            eventMiss.recordEvent(cpu_iid, tagged Invalid);
            stage5Ctrl.ready(cpu_iid, tuple3(local_state, tagged Invalid, ?));
        end
    endrule
    

    (* conservative_implicit_conditions *)
    rule stage4_STALL (stage4Stall matches tagged Valid {.cpu_iid,
                                                         .req,
                                                         .entry,
                                                         .ls});
        let local_state = ls;

        //
        // All events here will use the low bit to indicate whether the operation
        // is a load (0) or a store (1).  The remainer of the event data is
        // whatever fits from the low bits of the PA.
        //
        Maybe#(EVENT_PARAM) evt_hit = tagged Invalid;
        Maybe#(EVENT_PARAM) evt_miss = tagged Invalid;
        Maybe#(CACHE_PROTOCOL_MSG) new_miss_tok_req = tagged Invalid;

        //
        // Is the line already in the cache?
        //
        if (entry.state matches tagged Valid .state)
        begin
            // Yes:  hit
            if (cacheMsg_IsReqStore(req))
            begin
                if (!local_state.writePortUsed)
                begin
                    // We're writeback, so we don't need the memQ.
                    // Note that we don't need to do an eviction check since
                    // we hit, so we'll just overwrite the existing value.
                    // In other words, the writes will be coalesced and only
                    // one writeback to memory will occur.
                    local_state.writePortUsed = True;
                    local_state.writePortIdx = entry.idx;
                    local_state.writePortData = initCacheEntryState(req.linePAddr,
                                                                    True,
                                                                    ?);

                    // No response to a store. Don't change the coreQData in
                    // case there was a fill.
                    statWriteHit.incr(cpu_iid);
                    evt_hit = tagged Valid resize({ req.linePAddr, 1'b1 });
                    debugLog.record(cpu_iid, $format("3: STORE HIT"));
                    reqFromCore.doDeq(cpu_iid);
                end
                else
                begin
                    // The store must retry because a fill happened and the
                    // cache's write port is busy.
                    statWriteRetry.incr(cpu_iid);
                    debugLog.record(cpu_iid, $format("3: STORE HIT RETRY"));
                    reqFromCore.noDeq(cpu_iid);
                end
            end
            else if (local_state.coreQNotFull && ! local_state.coreQUsed)
            begin
                // A load hit, so give the data back. We won't need the
                // memory queue.
                local_state.coreQData = cacheMsg_RspLoad(req.linePAddr, req.opaque);
                local_state.coreQUsed = True;
                statReadHit.incr(cpu_iid);
                evt_hit = tagged Valid resize({ req.linePAddr, 1'b0 });
                debugLog.record(cpu_iid, $format("3: LOAD HIT"));
                reqFromCore.doDeq(cpu_iid);
            end
            else
            begin
                // A load hit, but the port is already in use, or the queue
                // is full, so retry.
                statReadRetry.incr(cpu_iid);
                debugLog.record(cpu_iid, $format("3: LOAD HIT RETRY"));
                reqFromCore.noDeq(cpu_iid);
            end
        end
        else
        begin
            //
            // Miss path.
            //
            if (entry.state matches tagged Blocked)
            begin
                // The request must stall because no line can currently be
                // evicted.
                statReadRetry.incr(cpu_iid);
                debugLog.record(cpu_iid, $format("3: EVICT BLOCKED RETRY"));
                reqFromCore.noDeq(cpu_iid);
            end
            else if (cacheMsg_IsReqStore(req))
            begin
                if (outstandingMisses.canAllocateStore(cpu_iid) &&
                    memQAvailable(local_state))
                begin
                    // Allocate the next miss ID.
                    new_miss_tok_req = tagged Valid req;
                    outstandingMisses.allocateStoreReq(cpu_iid);

                    // Record that we are using the memory queue.
                    local_state.memQUsed = True;

                    // A miss, so no response. (Don't change the response in case there's an existing fill)
                    //statWriteMiss.incr(cpu_iid);
                    evt_miss = tagged Valid resize({ req.linePAddr, 1'b1 });
                    debugLog.record(cpu_iid, $format("3: STORE MISS: ") + fshow(req));
                    reqFromCore.doDeq(cpu_iid);
                end
                else
                begin
                    // The request must stall.
                    statWriteRetry.incr(cpu_iid);
                    debugLog.record(cpu_iid, $format("3: STORE MISS RETRY"));
                    reqFromCore.noDeq(cpu_iid);
                end
            end
            else
            begin
                // A load miss. But do we have a free missID to track the fill?
                // And is the memQ not full and free for us to use?
                if (outstandingMisses.canAllocateLoad(cpu_iid) &&
                    memQAvailable(local_state))
                begin
                    // Allocate the next miss ID.
                    new_miss_tok_req = tagged Valid req;
                    outstandingMisses.allocateLoadReq(cpu_iid, req.linePAddr);

                    // Record that we are using the memory queue.
                    local_state.memQUsed = True;

                    // A miss, so no response. (Don't change the response in case
                    // there's an existing fill.)
                    statReadMiss.incr(cpu_iid);
                    evt_miss = tagged Valid resize({ req.linePAddr, 1'b0 });
                    debugLog.record(cpu_iid, $format("3: LOAD MISS: ") + fshow(req));
                    reqFromCore.doDeq(cpu_iid);
                end
                else
                begin
                    // The request must stall.
                    statReadRetry.incr(cpu_iid);
                    debugLog.record(cpu_iid, $format("3: LOAD MISS RETRY"));
                    reqFromCore.noDeq(cpu_iid);
                end
            end // cache load miss
        end
        
        eventHit.recordEvent(cpu_iid, evt_hit);
        eventMiss.recordEvent(cpu_iid, evt_miss);

        stage4Stall <= tagged Invalid;
        stage5Ctrl.ready(cpu_iid, tuple3(local_state, new_miss_tok_req, entry.idx));
    endrule
    

    rule stage5_end (True);
        match {.cpu_iid, {.local_state,
                          .new_miss_tok_req,
                          .fill_idx}} <- stage5Ctrl.nextReadyInstance();

        if (new_miss_tok_req matches tagged Valid .req)
        begin
            if (cacheMsg_IsReqStore(req))
            begin
                let miss_tok <- outstandingMisses.allocateStoreRsp(cpu_iid);

                // Record the cache index to which the fill will be written
                opaquesPool.write(cpu_iid, missTokIndex(miss_tok),
                                  tuple2(?, fill_idx));

                // Use the opaque bits to store the miss token.
                // Note that we use a load to simulate getting exclusive access.
                let mem_req = cacheMsg_ReqLoad(req.linePAddr,
                                               updateMemOpaque(req.opaque, miss_tok));
                local_state.memQData = mem_req;

                debugLog.record(cpu_iid, $format("4: STORE MISS: %0d, ", miss_tok.index) + fshow(req));
            end
            else
            begin
                let miss_tok <- outstandingMisses.allocateLoadRsp(cpu_iid);

                // Record the state of the outstanding fill, including the
                // L1 opaque.
                opaquesPool.write(cpu_iid, missTokIndex(miss_tok),
                                  tuple2(fromMemOpaque(req.opaque), fill_idx));

                // Use the opaque bits to store the miss token.
                let mem_req = cacheMsg_ReqLoad(req.linePAddr,
                                               updateMemOpaque(req.opaque, miss_tok));
                local_state.memQData = mem_req;

                debugLog.record(cpu_iid, $format("4: LOAD MISS: %0d, ", miss_tok.index) + fshow(req));
            end
        end

        // Take care of the memory queue.
        if (local_state.memQUsed)
        begin
            let req = local_state.memQData;
            let mreq = MEMORY_REQ { linePAddr: req.linePAddr,
                                    opaque: req.opaque,
                                    isStore: cacheMsg_IsReqStore(req) };

            reqToUncore.doEnq(cpu_iid, mreq);
        end
        else
        begin
            reqToUncore.noEnq(cpu_iid);
        end

        // Take care of the cache update.
        if (local_state.writePortUsed)
        begin
            if (! local_state.writePortData.dirty)
            begin
                // Fill -- must be an allocation
                l2Alg.allocate(cpu_iid,
                               local_state.writePortIdx,
                               local_state.writePortData,
                               CACHE_ALLOC_FILL);
            end
            else
            begin
                // Store.  In this controller, the line was already present.
                l2Alg.update(cpu_iid,
                             local_state.writePortIdx,
                             local_state.writePortData);
            end
        end

        // Take care of CPU rsp
        if (local_state.coreQUsed)
        begin
            rspToCore.doEnq(cpu_iid, local_state.coreQData);
        end
        else
        begin
            rspToCore.noEnq(cpu_iid);
        end

        // End of model cycle. (Path 1)
        debugLog.record(cpu_iid, $format("4: END CYCLE"));
        localCtrl.endModelCycle(cpu_iid, 1); 
    endrule
endmodule
