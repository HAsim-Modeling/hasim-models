
import hasim_common::*;
import hasim_modellib::*;

typedef NUM_CONTEXTS NUM_CPUS;
typedef INSTANCE_ID#(NUM_CPUS) CPU_INSTANCE_ID;

