`include "hasim_common.bsh"

module [HASIM_MODULE] mkSharedCache();
    return ?;
endmodule
