`include "asim/provides/hasim_common.bsh"

module [HASIM_MODULE] mkLastLevelCache();
endmodule
